library verilog;
use verilog.vl_types.all;
entity NivelRT_vlg_vec_tst is
end NivelRT_vlg_vec_tst;
